
`include "SRAM_wrapper.sv"
`include "CPU_wrapper.sv"
`include "./AXI/AXI.sv"
`include "DRAM_wrapper.sv"
`include "DMA_wrapper.sv"
`include "ROM_wrapper.sv"
`include "WDT_wrapper.sv"

module top (
	input clk,
	input rst,
	input clk2,
	input rst2, 
	input [31:0] DRAM_Q,
	input DRAM_valid,
	input [31:0] ROM_out,
	// DRAM
	output logic DRAM_CSn,
	output logic [3:0] DRAM_WEn,
	output logic DRAM_RASn,
	output logic DRAM_CASn,
	output logic [10:0] DRAM_A,
	output logic [31:0] DRAM_D,
	
	// ROM
	
	output logic ROM_read,
	output logic ROM_enable,
	output logic [11:0] ROM_address
);


logic [`AXI_ID_BITS-1:0] AWID_M0, AWID_M1, AWID_dma;
logic [`AXI_ADDR_BITS-1:0] AWADDR_M0, AWADDR_M1, AWADDR_dma;
logic [`AXI_LEN_BITS-1:0] AWLEN_M0, AWLEN_M1, AWLEN_dma;
logic [`AXI_SIZE_BITS-1:0] AWSIZE_M0, AWSIZE_M1, AWSIZE_dma;
logic [1:0] AWBURST_M0, AWBURST_M1, AWBURST_dma;
logic AWVALID_M0, AWVALID_M1, AWVALID_dma;
logic AWREADY_M0, AWREADY_M1, AWREADY_dma;
logic [`AXI_DATA_BITS-1:0] WDATA_M0, WDATA_M1, WDATA_dma;
logic [`AXI_STRB_BITS-1:0] WSTRB_M0, WSTRB_M1, WSTRB_dma;
logic WLAST_M0, WLAST_M1, WLAST_dma;
logic WVALID_M0, WVALID_M1, WVALID_dma;
logic WREADY_M0, WREADY_M1, WREADY_dma;
logic [`AXI_ID_BITS-1:0] BID_M0, BID_M1, BID_dma;
logic [1:0] BRESP_M0, BRESP_M1, BRESP_dma;
logic BVALID_M0, BVALID_M1, BVALID_dma;
logic BREADY_M0, BREADY_M1, BREADY_dma;
logic [`AXI_ID_BITS-1:0] ARID_M0, ARID_M1, ARID_dma;
logic [`AXI_ADDR_BITS-1:0] ARADDR_M0, ARADDR_M1, ARADDR_dma;
logic [`AXI_LEN_BITS-1:0] ARLEN_M0, ARLEN_M1, ARLEN_dma;
logic [`AXI_SIZE_BITS-1:0] ARSIZE_M0, ARSIZE_M1, ARSIZE_dma;
logic [1:0] ARBURST_M0, ARBURST_M1, ARBURST_dma;
logic ARVALID_M0, ARVALID_M1, ARVALID_dma;
logic ARREADY_M0, ARREADY_M1, ARREADY_dma;
logic [`AXI_ID_BITS-1:0] RID_M0, RID_M1, RID_dma;
logic [`AXI_DATA_BITS-1:0] RDATA_M0, RDATA_M1, RDATA_dma;
logic [1:0] RRESP_M0, RRESP_M1, RRESP_dma;
logic RLAST_M0, RLAST_M1, RLAST_dma;
logic RVALID_M0, RVALID_M1, RVALID_dma;
logic RREADY_M0, RREADY_M1, RREADY_dma;

logic [`AXI_IDS_BITS-1:0] ARID_S0;
logic [`AXI_ADDR_BITS-1:0] ARADDR_S0;
logic [`AXI_LEN_BITS-1:0] ARLEN_S0;
logic [`AXI_SIZE_BITS-1:0] ARSIZE_S0;
logic [1:0] ARBURST_S0;
logic ARVALID_S0;
logic ARREADY_S0;
logic [`AXI_IDS_BITS-1:0] RID_S0;
logic [`AXI_DATA_BITS-1:0] RDATA_S0;
logic [1:0] RRESP_S0;
logic RLAST_S0;
logic RVALID_S0;
logic RREADY_S0;
logic [`AXI_IDS_BITS-1:0] ARID_S1, ARID_S2, ARID_S3, ARID_S4, ARID_S5;
logic [`AXI_ADDR_BITS-1:0] ARADDR_S1, ARADDR_S2, ARADDR_S3, ARADDR_S4, ARADDR_S5;
logic [`AXI_LEN_BITS-1:0] ARLEN_S1, ARLEN_S2, ARLEN_S3, ARLEN_S4, ARLEN_S5;
logic [`AXI_SIZE_BITS-1:0] ARSIZE_S1, ARSIZE_S2, ARSIZE_S3, ARSIZE_S4, ARSIZE_S5;
logic [1:0] ARBURST_S1, ARBURST_S2, ARBURST_S3, ARBURST_S4, ARBURST_S5;
logic ARVALID_S1, ARVALID_S2, ARVALID_S3, ARVALID_S4, ARVALID_S5;
logic ARREADY_S1, ARREADY_S2, ARREADY_S3, ARREADY_S4, ARREADY_S5;
logic [`AXI_IDS_BITS-1:0] RID_S1, RID_S2, RID_S3, RID_S4, RID_S5;
logic [`AXI_DATA_BITS-1:0] RDATA_S1, RDATA_S2, RDATA_S3, RDATA_S4, RDATA_S5;
logic [1:0] RRESP_S1, RRESP_S2, RRESP_S3, RRESP_S4, RRESP_S5;
logic RLAST_S1, RLAST_S2, RLAST_S3, RLAST_S4, RLAST_S5;
logic RVALID_S1, RVALID_S2, RVALID_S3, RVALID_S4, RVALID_S5;
logic RREADY_S1, RREADY_S2, RREADY_S3, RREADY_S4, RREADY_S5;
logic [`AXI_IDS_BITS-1:0] AWID_S1, AWID_S2, AWID_S3, AWID_S4, AWID_S5;
logic [`AXI_ADDR_BITS-1:0] AWADDR_S1, AWADDR_S2, AWADDR_S3, AWADDR_S4, AWADDR_S5;
logic [`AXI_LEN_BITS-1:0] AWLEN_S1, AWLEN_S2, AWLEN_S3, AWLEN_S4, AWLEN_S5;
logic [`AXI_SIZE_BITS-1:0] AWSIZE_S1, AWSIZE_S2, AWSIZE_S3, AWSIZE_S4, AWSIZE_S5;
logic [1:0] AWBURST_S1, AWBURST_S2, AWBURST_S3, AWBURST_S4, AWBURST_S5;
logic AWVALID_S1, AWVALID_S2, AWVALID_S3, AWVALID_S4, AWVALID_S5;
logic AWREADY_S1, AWREADY_S2, AWREADY_S3, AWREADY_S4, AWREADY_S5;
logic [`AXI_DATA_BITS-1:0] WDATA_S1, WDATA_S2, WDATA_S3, WDATA_S4, WDATA_S5;
logic [`AXI_STRB_BITS-1:0] WSTRB_S1, WSTRB_S2, WSTRB_S3, WSTRB_S4, WSTRB_S5;
logic WLAST_S1, WLAST_S2, WLAST_S3, WLAST_S4, WLAST_S5;
logic WVALID_S1, WVALID_S2, WVALID_S3, WVALID_S4, WVALID_S5;
logic WREADY_S1, WREADY_S2, WREADY_S3, WREADY_S4, WREADY_S5;
logic [`AXI_IDS_BITS-1:0] BID_S1, BID_S2, BID_S3, BID_S4, BID_S5;
logic [1:0] BRESP_S1, BRESP_S2, BRESP_S3, BRESP_S4, BRESP_S5;
logic BVALID_S1, BVALID_S2, BVALID_S3, BVALID_S4, BVALID_S5;
logic BREADY_S1, BREADY_S2, BREADY_S3, BREADY_S4, BREADY_S5;
logic interrupt_dma, interrupt_time;
logic DMA_interrupt;

	

CPU_wrapper cpu(
	//input
	.ACLK(clk),
	.ARESETn(~rst),
	//WRITE ADDRESS1
	.AWID_M1(AWID_M1),
	.AWADDR_M1(AWADDR_M1),
	.AWLEN_M1(AWLEN_M1),
	.AWSIZE_M1(AWSIZE_M1),
	.AWBURST_M1(AWBURST_M1),
	.AWVALID_M1(AWVALID_M1),
	.AWREADY_M1(AWREADY_M1), //input
	//WRITE DATA1
	.WDATA_M1(WDATA_M1),
	.WSTRB_M1(WSTRB_M1),
	.WLAST_M1(WLAST_M1),
	.WVALID_M1(WVALID_M1),
	.WREADY_M1(WREADY_M1), //OUTPUT
	//WRITE RESPONSE1
	.BID_M1(BID_M1),
	.BRESP_M1(BRESP_M1),
	.BVALID_M1(BVALID_M1),
	.BREADY_M1(BREADY_M1), //OUTPUT
	//READ ADDRESS0
	.ARID_M0(ARID_M0),
	.ARADDR_M0(ARADDR_M0),
	.ARLEN_M0(ARLEN_M0),
	.ARSIZE_M0(ARSIZE_M0),
	.ARBURST_M0(ARBURST_M0),
	.ARVALID_M0(ARVALID_M0),
	.ARREADY_M0(ARREADY_M0), //INPUT
	//READ DATA0
	.RID_M0(RID_M0),
	.RDATA_M0(RDATA_M0),
	.RRESP_M0(RRESP_M0),
	.RLAST_M0(RLAST_M0),
	.RVALID_M0(RVALID_M0),
	.RREADY_M0(RREADY_M0), //OUTPUT
	//READ ADDRESS1
 	.ARID_M1(ARID_M1),
	.ARADDR_M1(ARADDR_M1),
	.ARLEN_M1(ARLEN_M1),
	.ARSIZE_M1(ARSIZE_M1),
	.ARBURST_M1(ARBURST_M1),
	.ARVALID_M1(ARVALID_M1),
	.ARREADY_M1(ARREADY_M1), //INPUT
	//READ DATA1
	.RID_M1(RID_M1),
	.RDATA_M1(RDATA_M1),
	.RRESP_M1(RRESP_M1),
	.RLAST_M1(RLAST_M1),
	.RVALID_M1(RVALID_M1),
	.RREADY_M1(RREADY_M1), //OUTPUT
	//interupt
	.interrupt_dma(DMA_interrupt),
	.interrupt_time(interrupt_time)
);

DMA_wrapper DMA(
	.ACLK(clk),
	.ARESETn(~rst),

	//WRITE ADDRESS1
	.AWID_dma(AWID_dma),
	.AWADDR_dma(AWADDR_dma),
	.AWLEN_dma(AWLEN_dma),
	.AWSIZE_dma(AWSIZE_dma),
	.AWBURST_dma(AWBURST_dma),
	.AWVALID_dma(AWVALID_dma),
	.AWREADY_dma(AWREADY_dma),
	
	//WRITE DATA1
	.WDATA_dma(WDATA_dma),
	.WSTRB_dma(WSTRB_dma),
	.WLAST_dma(WLAST_dma),
	.WVALID_dma(WVALID_dma),
	.WREADY_dma(WREADY_dma),
	
	//WRITE RESPONSE1
	.BID_dma(BID_dma),
	.BRESP_dma(BRESP_dma),
	.BVALID_dma(BVALID_dma),
	.BREADY_dma(BREADY_dma),

	//READ ADDRESS0
	.ARID_dma(ARID_dma),
	.ARADDR_dma(ARADDR_dma),
	.ARLEN_dma(ARLEN_dma),
	.ARSIZE_dma(ARSIZE_dma),
	.ARBURST_dma(ARBURST_dma),
	.ARVALID_dma(ARVALID_dma),
	.ARREADY_dma(ARREADY_dma),
	
	//READ DATA0
	.RID_dma(RID_dma),
	.RDATA_dma(RDATA_dma),
	.RRESP_dma(RRESP_dma),
	.RLAST_dma(RLAST_dma),
	.RVALID_dma(RVALID_dma),
	.RREADY_dma(RREADY_dma),

	//SLAVE INTERFACE FOR MASTERS
	
	//WRITE ADDRESS
	.AWID_S(AWID_S3),
	.AWADDR_S(AWADDR_S3),
	.AWLEN_S(AWLEN_S3),
	.AWSIZE_S(AWSIZE_S3),
	.AWBURST_S(AWBURST_S3),
	.AWVALID_S(AWVALID_S3),
	.AWREADY_S(AWREADY_S3),
	
	//WRITE DATA
	.WDATA_S(WDATA_S3),
	.WSTRB_S(WSTRB_S3),
	.WLAST_S(WLAST_S3),
	.WVALID_S(WVALID_S3),
	.WREADY_S(WREADY_S3),
	
	//WRITE RESPONSE
	.BID_S(BID_S3),
	.BRESP_S(BRESP_S3),
	.BVALID_S(BVALID_S3),
	.BREADY_S(BREADY_S3),

	//READ ADDRESS0
	.ARID_S(ARID_S3),
	.ARADDR_S(ARADDR_S3),
	.ARLEN_S(ARLEN_S3),
	.ARSIZE_S(ARSIZE_S3),
	.ARBURST_S(ARBURST_S3),
	.ARVALID_S(ARVALID_S3),
	.ARREADY_S(ARREADY_S3),
	
	//READ DATA0
	.RID_S(RID_S3),
	.RDATA_S(RDATA_S3),
	.RRESP_S(RRESP_S3),
	.RLAST_S(RLAST_S3),
	.RVALID_S(RVALID_S3),
	.RREADY_S(RREADY_S3),
	//
	.DMA_interrupt(DMA_interrupt)
	
);

AXI axi(
	.ACLK(clk),
	.ARESETn(~rst),
	//slave
	//read address 0
	.ARID_M0(ARID_M0),
	.ARADDR_M0(ARADDR_M0),
	.ARLEN_M0(ARLEN_M0),
	.ARSIZE_M0(ARSIZE_M0),
	.ARBURST_M0(ARBURST_M0),
	.ARVALID_M0(ARVALID_M0),
	.ARREADY_M0(ARREADY_M0),
	//READ DATA0
	.RID_M0(RID_M0),
	.RDATA_M0(RDATA_M0),
	.RRESP_M0(RRESP_M0),
	.RLAST_M0(RLAST_M0),
	.RVALID_M0(RVALID_M0),
	.RREADY_M0(RREADY_M0),
	//READ ADDRESS1
	.ARID_M1(ARID_M1),
	.ARADDR_M1(ARADDR_M1),
	.ARLEN_M1(ARLEN_M1),
	.ARSIZE_M1(ARSIZE_M1),
	.ARBURST_M1(ARBURST_M1),
	.ARVALID_M1(ARVALID_M1),
	.ARREADY_M1(ARREADY_M1),
	//READ DATA1
	.RID_M1(RID_M1),
	.RDATA_M1(RDATA_M1),
	.RRESP_M1(RRESP_M1),
	.RLAST_M1(RLAST_M1),
	.RVALID_M1(RVALID_M1),
	.RREADY_M1(RREADY_M1),
	//WRITE ADDRESS
	.AWID_M1(AWID_M1),
	.AWADDR_M1(AWADDR_M1),
	.AWLEN_M1(AWLEN_M1),
	.AWSIZE_M1(AWSIZE_M1),
	.AWBURST_M1(AWBURST_M1),
	.AWVALID_M1(AWVALID_M1),
	.AWREADY_M1(AWREADY_M1),
	//WRITE DATA
	.WDATA_M1(WDATA_M1),
	.WSTRB_M1(WSTRB_M1),
	.WLAST_M1(WLAST_M1),
	.WVALID_M1(WVALID_M1),
	.WREADY_M1(WREADY_M1),
	//WRITE RESPONSE
	.BID_M1(BID_M1),
	.BRESP_M1(BRESP_M1),
	.BVALID_M1(BVALID_M1),
	.BREADY_M1(BREADY_M1),

	//WRITE ADDRESS dma
	.AWID_dma(AWID_dma),
	.AWADDR_dma(AWADDR_dma),
	.AWLEN_dma(AWLEN_dma),
	.AWSIZE_dma(AWSIZE_dma),
	.AWBURST_dma(AWBURST_dma),
	.AWVALID_dma(AWVALID_dma),
	.AWREADY_dma(AWREADY_dma),
	
	//WRITE DATA dma
	.WDATA_dma(WDATA_dma),
	.WSTRB_dma(WSTRB_dma),
	.WLAST_dma(WLAST_dma),
	.WVALID_dma(WVALID_dma),
	.WREADY_dma(WREADY_dma),
	
	//WRITE RESPONSE dma
	.BID_dma(BID_dma),
	.BRESP_dma(BRESP_dma),
	.BVALID_dma(BVALID_dma),
	.BREADY_dma(BREADY_dma),

	//READ ADDRESS0
	.ARID_dma(ARID_dma),
	.ARADDR_dma(ARADDR_dma),
	.ARLEN_dma(ARLEN_dma),
	.ARSIZE_dma(ARSIZE_dma),
	.ARBURST_dma(ARBURST_dma),
	.ARVALID_dma(ARVALID_dma),
	.ARREADY_dma(ARREADY_dma),
	
	//READ DATA0
	.RID_dma(RID_dma),
	.RDATA_dma(RDATA_dma),
	.RRESP_dma(RRESP_dma),
	.RLAST_dma(RLAST_dma),
	.RVALID_dma(RVALID_dma),
	.RREADY_dma(RREADY_dma),

	//MASTER
	//READ ADDRESS 0
	.ARID_S0(ARID_S0),
	.ARADDR_S0(ARADDR_S0),
	.ARLEN_S0(ARLEN_S0),
	.ARSIZE_S0(ARSIZE_S0),
	.ARBURST_S0(ARBURST_S0),
	.ARVALID_S0(ARVALID_S0),
	.ARREADY_S0(ARREADY_S0),
	//READ DATA0
	.RID_S0(RID_S0),
	.RDATA_S0(RDATA_S0),
	.RRESP_S0(RRESP_S0),
	.RLAST_S0(RLAST_S0),
	.RVALID_S0(RVALID_S0),
	.RREADY_S0(RREADY_S0),
	//READ ADDRESS1
	.ARID_S1(ARID_S1),
	.ARADDR_S1(ARADDR_S1),
	.ARLEN_S1(ARLEN_S1),
	.ARSIZE_S1(ARSIZE_S1),
	.ARBURST_S1(ARBURST_S1),
	.ARVALID_S1(ARVALID_S1),
	.ARREADY_S1(ARREADY_S1),
	//READ DATA1
	.RID_S1(RID_S1),
	.RDATA_S1(RDATA_S1),
	.RRESP_S1(RRESP_S1),
	.RLAST_S1(RLAST_S1),
	.RVALID_S1(RVALID_S1),
	.RREADY_S1(RREADY_S1),
	//READ ADDRESS3
	.ARID_S2(ARID_S2),
	.ARADDR_S2(ARADDR_S2),
	.ARLEN_S2(ARLEN_S2),
	.ARSIZE_S2(ARSIZE_S2),
	.ARBURST_S2(ARBURST_S2),
	.ARVALID_S2(ARVALID_S2),
	.ARREADY_S2(ARREADY_S2),
	//READ DATA3
	.RID_S2(RID_S2),
	.RDATA_S2(RDATA_S2),
	.RRESP_S2(RRESP_S2),
	.RLAST_S2(RLAST_S2),
	.RVALID_S2(RVALID_S2),
	.RREADY_S2(RREADY_S2),
	//READ ADDRESS3
	.ARID_S3(ARID_S3),
	.ARADDR_S3(ARADDR_S3),
	.ARLEN_S3(ARLEN_S3),
	.ARSIZE_S3(ARSIZE_S3),
	.ARBURST_S3(ARBURST_S3),
	.ARVALID_S3(ARVALID_S3),
	.ARREADY_S3(ARREADY_S3),
	//READ DATA3
	.RID_S3(RID_S3),
	.RDATA_S3(RDATA_S3),
	.RRESP_S3(RRESP_S3),
	.RLAST_S3(RLAST_S3),
	.RVALID_S3(RVALID_S3),
	.RREADY_S3(RREADY_S3),
	
	//READ ADDRESS5
	.ARID_S5(ARID_S5),
	.ARADDR_S5(ARADDR_S5),
	.ARLEN_S5(ARLEN_S5),
	.ARSIZE_S5(ARSIZE_S5),
	.ARBURST_S5(ARBURST_S5),
	.ARVALID_S5(ARVALID_S5),
	.ARREADY_S5(ARREADY_S5),
	//READ DATA5
	.RID_S5(RID_S5),
	.RDATA_S5(RDATA_S5),
	.RRESP_S5(RRESP_S5),
	.RLAST_S5(RLAST_S5),
	.RVALID_S5(RVALID_S5),
	.RREADY_S5(RREADY_S5),
	//WRITE ADDRESS0
	.AWID_S1(AWID_S1),
	.AWADDR_S1(AWADDR_S1),
	.AWLEN_S1(AWLEN_S1),
	.AWSIZE_S1(AWSIZE_S1),
	.AWBURST_S1(AWBURST_S1),
	.AWVALID_S1(AWVALID_S1),
	.AWREADY_S1(AWREADY_S1),
	//WRITE DATA0
	.WDATA_S1(WDATA_S1),
	.WSTRB_S1(WSTRB_S1),
	.WLAST_S1(WLAST_S1),
	.WVALID_S1(WVALID_S1),
	.WREADY_S1(WREADY_S1),
	//WRITE RESPONSE0
	.BID_S1(BID_S1),
	.BRESP_S1(BRESP_S1),
	.BVALID_S1(BVALID_S1),
	.BREADY_S1(BREADY_S1),
	//WRITE ADDRESS2
	.AWID_S2(AWID_S2),
	.AWADDR_S2(AWADDR_S2),
	.AWLEN_S2(AWLEN_S2),
	.AWSIZE_S2(AWSIZE_S2),
	.AWBURST_S2(AWBURST_S2),
	.AWVALID_S2(AWVALID_S2),
	.AWREADY_S2(AWREADY_S2),
	//WRITE DATA2
	.WDATA_S2(WDATA_S2),
	.WSTRB_S2(WSTRB_S2),	
	.WLAST_S2(WLAST_S2),
	.WVALID_S2(WVALID_S2),
	.WREADY_S2(WREADY_S2),
	.BID_S2(BID_S2),
	.BRESP_S2(BRESP_S2),
	.BVALID_S2(BVALID_S2),
	.BREADY_S2(BREADY_S2),
	//WRITE ADDRESS3
	.AWID_S3(AWID_S3),
	.AWADDR_S3(AWADDR_S3),
	.AWLEN_S3(AWLEN_S3),
	.AWSIZE_S3(AWSIZE_S3),
	.AWBURST_S3(AWBURST_S3),
	.AWVALID_S3(AWVALID_S3),
	.AWREADY_S3(AWREADY_S3),
	//WRITE DATA3
	.WDATA_S3(WDATA_S3),
	.WSTRB_S3(WSTRB_S3),	
	.WLAST_S3(WLAST_S3),
	.WVALID_S3(WVALID_S3),
	.WREADY_S3(WREADY_S3),
	.BID_S3(BID_S3),
	.BRESP_S3(BRESP_S3),
	.BVALID_S3(BVALID_S3),
	.BREADY_S3(BREADY_S3),
	//WRITE ADDRESS4
	.AWID_S4(AWID_S4),
	.AWADDR_S4(AWADDR_S4),
	.AWLEN_S4(AWLEN_S4),
	.AWSIZE_S4(AWSIZE_S4),
	.AWBURST_S4(AWBURST_S4),
	.AWVALID_S4(AWVALID_S4),
	.AWREADY_S4(AWREADY_S4),
	//WRITE DATA4
	.WDATA_S4(WDATA_S4),
	.WSTRB_S4(WSTRB_S4),	
	.WLAST_S4(WLAST_S4),
	.WVALID_S4(WVALID_S4),
	.WREADY_S4(WREADY_S4),
	.BID_S4(BID_S4),
	.BRESP_S4(BRESP_S4),
	.BVALID_S4(BVALID_S4),
	.BREADY_S4(BREADY_S4),
	//WRITE ADDRESS5
	.AWID_S5(AWID_S5),
	.AWADDR_S5(AWADDR_S5),
	.AWLEN_S5(AWLEN_S5),
	.AWSIZE_S5(AWSIZE_S5),
	.AWBURST_S5(AWBURST_S5),
	.AWVALID_S5(AWVALID_S5),
	.AWREADY_S5(AWREADY_S5),
	//WRITE DATA5
	.WDATA_S5(WDATA_S5),
	.WSTRB_S5(WSTRB_S5),	
	.WLAST_S5(WLAST_S5),
	.WVALID_S5(WVALID_S5),
	.WREADY_S5(WREADY_S5),
	.BID_S5(BID_S5),
	.BRESP_S5(BRESP_S5),
	.BVALID_S5(BVALID_S5),
	.BREADY_S5(BREADY_S5)
);


SRAM_wrapper IM1(
	.ACLK(clk),
	.ARESETn(~rst),
	//WRITE ADDRESS
	.AWID_S(AWID_S1),
	.AWADDR_S(AWADDR_S1),
	.AWLEN_S(AWLEN_S1),
	.AWSIZE_S(AWSIZE_S1),
	.AWBURST_S(AWBURST_S1),
	.AWVALID_S(AWVALID_S1),	
	.AWREADY_S(AWREADY_S1), //output
	//WRITE DATA
	.WDATA_S(WDATA_S1),	
	.WSTRB_S(WSTRB_S1),
	.WLAST_S(WLAST_S1),
	.WVALID_S(WVALID_S1),
	.WREADY_S(WREADY_S1),  //output
	//WRITE RESPONSE
	.BID_S(BID_S1),
	.BRESP_S(BRESP_S1),
	.BVALID_S(BVALID_S1),	
	.BREADY_S(BREADY_S1),  //input
	//READ ADDRESS0
	.ARID_S(ARID_S1),
	.ARADDR_S(ARADDR_S1),
	.ARLEN_S(ARLEN_S1),
	.ARSIZE_S(ARSIZE_S1),
	.ARBURST_S(ARBURST_S1),
	.ARVALID_S(ARVALID_S1),
	.ARREADY_S(ARREADY_S1),  //output
	//READ DATA0
	.RID_S(RID_S1),	
	.RDATA_S(RDATA_S1),
	.RRESP_S(RRESP_S1),
	.RLAST_S(RLAST_S1),
	.RVALID_S(RVALID_S1),
	.RREADY_S(RREADY_S1)  //input
);

SRAM_wrapper DM1(
	.ACLK(clk),
	.ARESETn(~rst),
	//WRITE ADDRESS1
	.AWID_S(AWID_S2),
	.AWADDR_S(AWADDR_S2),
	.AWLEN_S(AWLEN_S2),
	.AWSIZE_S(AWSIZE_S2),
	.AWBURST_S(AWBURST_S2),
	.AWVALID_S(AWVALID_S2),	
	.AWREADY_S(AWREADY_S2), //output
	//WRITE DATA1
	.WDATA_S(WDATA_S2),	
	.WSTRB_S(WSTRB_S2),
	.WLAST_S(WLAST_S2),
	.WVALID_S(WVALID_S2),
	.WREADY_S(WREADY_S2),  //output
	//WRITE RESPONSE1
	.BID_S(BID_S2),
	.BRESP_S(BRESP_S2),
	.BVALID_S(BVALID_S2),	
	.BREADY_S(BREADY_S2),  //input
	//READ ADDRESS1
	.ARID_S(ARID_S2),
	.ARADDR_S(ARADDR_S2),
	.ARLEN_S(ARLEN_S2),
	.ARSIZE_S(ARSIZE_S2),
	.ARBURST_S(ARBURST_S2),
	.ARVALID_S(ARVALID_S2),
	.ARREADY_S(ARREADY_S2),  //output
	//READ DATA1
	.RID_S(RID_S2),	
	.RDATA_S(RDATA_S2),
	.RRESP_S(RRESP_S2),
	.RLAST_S(RLAST_S2),
	.RVALID_S(RVALID_S2),
	.RREADY_S(RREADY_S2)  //input
);

DRAM_wrapper DRAM(
	.ACLK(clk),
	.ARESETn(~rst),
	//WRITE ADDRESS3
	.AWID_S(AWID_S5),
	.AWADDR_S(AWADDR_S5),
	.AWLEN_S(AWLEN_S5),
	.AWSIZE_S(AWSIZE_S5),
	.AWBURST_S(AWBURST_S5),
	.AWVALID_S(AWVALID_S5),	
	.AWREADY_S(AWREADY_S5), //output
	//WRITE DATA3
	.WDATA_S(WDATA_S5),	
	.WSTRB_S(WSTRB_S5),
	.WLAST_S(WLAST_S5),
	.WVALID_S(WVALID_S5),
	.WREADY_S(WREADY_S5),  //output
	//WRITE RESPONSE3
	.BID_S(BID_S5),
	.BRESP_S(BRESP_S5),
	.BVALID_S(BVALID_S5),	
	.BREADY_S(BREADY_S5),  //input
	//READ ADDRESS3
	.ARID_S(ARID_S5),
	.ARADDR_S(ARADDR_S5),
	.ARLEN_S(ARLEN_S5),
	.ARSIZE_S(ARSIZE_S5),
	.ARBURST_S(ARBURST_S5),
	.ARVALID_S(ARVALID_S5),
	.ARREADY_S(ARREADY_S5),  //output
	//READ DATA3
	.RID_S(RID_S5),	
	.RDATA_S(RDATA_S5),
	.RRESP_S(RRESP_S5),
	.RLAST_S(RLAST_S5),
	.RVALID_S(RVALID_S5),
	.RREADY_S(RREADY_S5),  //input
	.CSn(DRAM_CSn),
	.WEn(DRAM_WEn),
	.RASn(DRAM_RASn),
	.CASn(DRAM_CASn),
	.A(DRAM_A),
	.D(DRAM_D),
	.Q(DRAM_Q),
	.valid(DRAM_valid)
);

ROM_wrapper ROM(
	.ACLK(clk),
	.ARESETn(~rst),
	//READ ADDRESS3
	.ARID_S(ARID_S0),
	.ARADDR_S(ARADDR_S0),
	.ARLEN_S(ARLEN_S0),
	.ARSIZE_S(ARSIZE_S0),
	.ARBURST_S(ARBURST_S0),
	.ARVALID_S(ARVALID_S0),
	.ARREADY_S(ARREADY_S0),  //output
	//READ DATA3
	.RID_S(RID_S0),	
	.RDATA_S(RDATA_S0),
	.RRESP_S(RRESP_S0),
	.RLAST_S(RLAST_S0),
	.RVALID_S(RVALID_S0),
	.RREADY_S(RREADY_S0),  //input
	.ROM_out(ROM_out),	//input
	.ROM_read(ROM_read),
	.ROM_enable(ROM_enable),
	.ROM_address(ROM_address)
);

WDT_wrapper WDT(
	.ACLK(clk),
	.ACLK2(clk2),
	.ARESETn(~rst),
	.ARESETn2(~rst2),
	//WRITE ADDRESS1
	.AWID_S(AWID_S4),
	.AWADDR_S(AWADDR_S4),
	.AWLEN_S(AWLEN_S4),
	.AWSIZE_S(AWSIZE_S4),
	.AWBURST_S(AWBURST_S4),
	.AWVALID_S(AWVALID_S4),	
	.AWREADY_S(AWREADY_S4), //output
	//WRITE DATA1
	.WDATA_S(WDATA_S4),	
	.WSTRB_S(WSTRB_S4),
	.WLAST_S(WLAST_S4),
	.WVALID_S(WVALID_S4),
	.WREADY_S(WREADY_S4),  //output
	//WRITE RESPONSE1
	.BID_S(BID_S4),
	.BRESP_S(BRESP_S4),
	.BVALID_S(BVALID_S4),	
	.BREADY_S(BREADY_S4), //input

	.WTO(interrupt_time)
	
);



endmodule

