`define CPU_CYCLE     1.9 // 100Mhz
`define MAX           300000000 // 3000000
